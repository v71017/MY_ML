0.8476469207350941
1 4.0 4.908008 2.52006
-1 4.0 0.537667 0.888396
1 4.0 2.825219 1.979972
-1 4.0 1.833885 -1.14707
-1 4.0 -2.258847 -1.06887
-1 4.0 3.578397 1.370299
1 4.0 1.738005 -0.329867
1 4.0 0.249788 0.550903
